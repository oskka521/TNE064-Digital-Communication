library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity img_gen is
	Port ( 
			 clk         : in  STD_LOGIC;
			 x_control   : in  STD_LOGIC_VECTOR(9 downto 0);
			 y_control   : in  STD_LOGIC_VECTOR(9 downto 0);
			 rgb         : out STD_LOGIC_VECTOR(3 downto 0)
			 );
end img_gen;

architecture Behavioral of img_gen is
	

	constant 	Xpos:								integer:=280; --	640/2 - 80/2 = 280
	constant 	Ypos:								integer:=210; --  480/2 - 60/2 = 210
	constant 	bredd:							integer:=80;
	constant 	hojd:								integer:=60;
	signal 		refresh_tick:					std_logic;
	

	signal x,y:integer range 0 to 650;
	signal rgb_reg,rgb_next:std_logic_vector(3 downto 0);
	signal counter:integer;
	
	type rom_type is array (0 to 4800 -1) of std_logic_vector (3 downto 0);  
	signal rom : rom_type:= ("0001", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0001", "0011", "0011", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0001", "0001", "0001", "0001", "0001", "0000", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0000", "0000", "0001", "0001", "0001", "0010", "0100", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0010", "0001", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0000", "0001", "0001", "0001", "0010", "0011", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0101", "0110", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "1000", "0011", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0000", "0001", "0001", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0010", "0100", "0100", "0100", "0101", "0101", "0101", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "1010", "1001", "0100", "0001", "0001", "0001", "0001", "0001", "0000", "0000", "0001", "0001", "0001", "0001", "0001", "0001", "0000", "0001", "0010", "0011", "0100", "0100", "0101", "0101", "0101", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0100", "0101", "0101", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0100", "0101", "0101", "1010", "1010", "1010", "0110", "0001", "0001", "0001", "0001", "0000", "0000", "0001", "0001", "0001", "0010", "0001", "0001", "0001", "0001", "0001", "0010", "0011", "0101", "0101", "0101", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1001", "1000", "1000", "0111", "0110", "0111", "1000", "1000", "0110", "0110", "0101", "0101", "0101", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "1001", "1001", "1010", "1010", "0101", "0001", "0010", "0001", "0001", "0000", "0000", "0001", "0010", "0010", "0010", "0010", "0001", "0001", "0001", "0001", "0010", "0100", "0101", "0101", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "1000", "1000", "0111", "0111", "1000", "1000", "1000", "0111", "1000", "1010", "1100", "1001", "0111", "0111", "0110", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0110", "0110", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0111", "1001", "1001", "1001", "1010", "1010", "0101", "0001", "0010", "0001", "0000", "0001", "0001", "0010", "0010", "0010", "0010", "0010", "0001", "0001", "0001", "0001", "0001", "0100", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "1000", "1000", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1011", "1001", "0111", "0111", "0111", "0111", "0110", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0101", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0110", "0111", "1010", "1010", "1010", "1001", "1001", "1001", "0110", "0011", "0001", "0000", "0001", "0001", "0001", "0010", "0011", "0011", "0011", "0001", "0001", "0001", "0001", "0011", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0110", "0110", "0101", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "0110", "0001", "0000", "0001", "0001", "0010", "0011", "0011", "0011", "0100", "0010", "0010", "0010", "0001", "0011", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "1000", "1000", "1001", "1001", "1010", "1010", "1010", "1010", "1001", "1010", "1010", "1010", "1010", "1001", "1000", "1000", "1000", "1001", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0101", "0101", "0101", "0101", "0101", "0101", "0111", "1000", "1010", "1010", "1010", "1010", "1010", "1010", "1100", "1011", "0100", "0000", "0010", "0010", "0001", "0010", "0010", "0011", "0100", "0100", "0011", "0011", "0011", "0101", "0110", "0110", "0111", "0111", "0111", "0111", "1000", "1000", "1001", "1001", "1001", "1010", "1011", "1011", "1011", "1010", "1010", "1011", "1011", "1011", "1010", "1001", "1001", "1010", "1010", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0101", "0101", "0101", "0110", "0110", "0110", "1000", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1011", "1011", "1011", "1010", "0010", "0011", "0011", "0010", "0001", "0001", "0001", "0010", "0100", "0100", "0011", "0101", "0110", "0110", "0110", "0111", "0111", "1000", "1000", "1000", "1001", "1001", "1001", "1010", "1010", "1011", "1100", "1100", "1011", "1011", "1011", "1011", "1010", "1010", "1001", "1001", "1001", "1001", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0110", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "1010", "1001", "1000", "1010", "1010", "1010", "1010", "1010", "1010", "1011", "1011", "1011", "0111", "0010", "0011", "0011", "0010", "0001", "0001", "0001", "0011", "0101", "0101", "0101", "0110", "0110", "0111", "0111", "0111", "1000", "1000", "1001", "1001", "1010", "1010", "1010", "1011", "1100", "1101", "1101", "1100", "1101", "1100", "1011", "1011", "1010", "1010", "1010", "1001", "1001", "1000", "1000", "1001", "1000", "0111", "0111", "0111", "0111", "1000", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "1000", "1000", "0111", "0111", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "0100", "0011", "0100", "0011", "0010", "0010", "0001", "0011", "0100", "0101", "0110", "0110", "0110", "0111", "0111", "1000", "1000", "1000", "1001", "1010", "1010", "1011", "1011", "1100", "1100", "1110", "1110", "1110", "1110", "1101", "1100", "1011", "1011", "1011", "1010", "1001", "1001", "1001", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "1000", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1000", "1010", "1010", "1010", "1010", "1011", "1011", "1010", "1010", "1010", "1010", "1001", "0101", "0100", "0100", "0010", "0010", "0010", "0001", "0011", "0110", "0110", "0110", "0111", "0111", "0111", "1000", "1000", "1000", "1001", "1001", "1010", "1011", "1100", "1101", "1101", "1110", "1111", "1111", "1111", "1101", "1101", "1101", "1100", "1011", "1010", "1010", "1001", "1001", "1000", "1000", "1000", "1000", "1010", "1011", "1001", "1010", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "1000", "0111", "0111", "1001", "1001", "1001", "1010", "1010", "1010", "1011", "1011", "1010", "1010", "1010", "1010", "1001", "0101", "0100", "0011", "0010", "0011", "0010", "0010", "0100", "0110", "0110", "0111", "0111", "0111", "1000", "1000", "1000", "1001", "1001", "1010", "1011", "1100", "1101", "1111", "1111", "1111", "1111", "1111", "1111", "1110", "1101", "1100", "1011", "1010", "1010", "1001", "1001", "1001", "1000", "1000", "1001", "1100", "1011", "1001", "1010", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0110", "0110", "0110", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "0111", "1000", "1011", "1011", "1010", "1001", "1001", "1010", "1010", "1011", "1011", "1011", "1010", "1010", "1011", "1001", "0100", "0100", "0010", "0010", "0011", "0011", "0100", "0110", "0110", "0111", "0111", "1000", "1000", "1000", "1001", "1001", "1010", "1010", "1011", "1100", "1101", "1110", "1111", "1111", "1111", "1111", "1111", "1101", "1100", "1100", "1011", "1010", "1010", "1001", "1010", "1010", "1001", "1001", "1001", "1011", "1001", "1001", "1001", "1001", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1001", "1100", "1101", "1100", "1100", "1100", "1011", "1010", "1010", "1010", "1011", "1011", "1011", "1011", "1011", "1010", "0101", "0100", "0100", "0011", "0011", "0011", "0101", "0110", "0111", "0111", "0111", "1000", "1000", "1000", "1001", "1001", "1010", "1011", "1011", "1100", "1110", "1111", "1111", "1111", "1111", "1111", "1111", "1110", "1101", "1100", "1011", "1010", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1010", "1100", "1011", "1010", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1001", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1101", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1010", "0110", "0101", "0100", "0011", "0011", "0110", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1001", "1001", "1010", "1011", "1100", "1101", "1101", "1110", "1110", "1111", "1111", "1111", "1110", "1110", "1101", "1100", "1011", "1011", "1010", "1010", "1001", "1010", "1010", "1010", "1010", "1011", "1100", "1100", "1010", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1010", "1101", "1110", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1100", "1100", "1100", "1011", "1011", "1011", "1100", "1011", "1000", "0101", "0101", "0101", "0110", "0111", "0111", "0111", "0111", "1000", "1000", "1000", "1001", "1001", "1010", "1011", "1011", "1100", "1100", "1101", "1110", "1110", "1110", "1111", "1110", "1101", "1100", "1100", "1011", "1011", "1011", "1100", "1100", "1001", "1001", "1001", "1010", "1011", "1100", "1011", "1010", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "0111", "0111", "0111", "0111", "0111", "1000", "1011", "1101", "1110", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1100", "1011", "1100", "1110", "1101", "1001", "0110", "0110", "0110", "0110", "0111", "0111", "0111", "1000", "1000", "1001", "1001", "1010", "1010", "1010", "1011", "1011", "1100", "1101", "1110", "1101", "1101", "1110", "1101", "1100", "1100", "1011", "1011", "1100", "1111", "1110", "1101", "1010", "1010", "1100", "1011", "1011", "1100", "1010", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "0111", "1000", "1000", "1010", "1101", "1110", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1110", "1110", "1011", "0111", "0110", "0111", "0111", "0111", "0111", "1000", "1000", "1001", "1001", "1001", "1010", "1010", "1010", "1011", "1011", "1100", "1101", "1100", "1100", "1101", "1101", "1100", "1011", "1011", "1011", "1101", "1110", "1101", "1100", "1011", "1011", "1100", "1011", "1010", "1010", "1001", "1000", "1000", "1001", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1010", "1101", "1110", "1110", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1111", "1101", "1000", "0110", "0111", "0111", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1010", "1010", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1011", "1100", "1101", "1101", "1011", "1011", "1010", "1010", "1011", "1001", "1001", "1001", "1010", "1011", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1001", "1101", "1110", "1110", "1101", "1100", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1111", "1110", "1001", "0111", "0111", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1001", "1010", "1010", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1011", "1011", "1100", "1101", "1101", "1101", "1011", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1010", "1001", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1000", "1001", "1010", "1101", "1110", "1110", "1110", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1111", "1110", "1011", "0111", "0111", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1010", "1010", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1110", "1101", "1100", "1010", "1101", "1011", "1001", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1000", "1000", "1001", "1001", "1001", "1000", "1000", "1001", "1001", "1010", "1101", "1110", "1110", "1101", "1101", "1101", "1101", "1110", "1101", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1111", "1111", "1100", "1001", "1000", "1000", "1000", "1000", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1011", "1011", "1011", "1011", "1011", "1110", "1101", "1101", "1100", "1011", "1011", "1010", "1010", "1011", "1010", "1001", "1010", "1001", "1001", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1011", "1110", "1110", "1110", "1100", "1100", "1101", "1101", "1110", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1111", "1110", "1110", "1100", "1001", "1000", "1000", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1011", "1100", "1100", "1011", "1011", "1010", "1011", "1011", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1011", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1001", "1010", "1100", "1110", "1110", "1110", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1100", "1100", "1100", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1110", "1110", "1110", "1110", "1111", "1110", "1110", "1110", "1100", "1001", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1011", "1100", "1011", "1100", "1100", "1011", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1010", "1011", "1011", "1010", "1010", "1010", "1010", "1010", "1001", "1001", "1001", "1001", "1011", "1110", "1110", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1111", "1110", "1110", "1110", "1100", "1001", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1011", "1011", "1011", "1101", "1100", "1011", "1010", "1010", "1010", "1011", "1010", "1001", "1010", "0111", "0100", "0110", "1011", "1100", "1101", "1101", "1010", "1001", "1010", "1010", "1011", "1110", "1110", "1101", "1101", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1101", "1101", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1110", "1110", "1101", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1111", "1111", "1111", "1110", "1100", "1010", "1010", "1001", "1001", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1011", "1011", "1011", "1011", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "0011", "0001", "0001", "1011", "1111", "1111", "1101", "1010", "1010", "1010", "1011", "1101", "1110", "1101", "1110", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1101", "1110", "1110", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1110", "1101", "1100", "1011", "1010", "1010", "1010", "1010", "1010", "1011", "1011", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1011", "1001", "0100", "0010", "0010", "0010", "1011", "1111", "1101", "1011", "1010", "1010", "1011", "1100", "1100", "1100", "1101", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1101", "1100", "1011", "1001", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "1010", "0101", "0010", "0001", "0010", "0010", "0111", "1101", "1011", "1011", "1011", "1100", "1100", "1011", "1011", "1101", "1110", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1110", "1110", "1101", "1101", "1011", "1100", "1101", "1100", "1100", "1101", "1001", "0011", "0011", "0001", "0001", "0001", "0001", "0101", "1011", "1100", "1011", "1100", "1011", "1101", "1110", "1110", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1100", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1111", "1111", "1110", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1110", "0111", "0100", "0011", "0010", "0010", "0010", "0001", "0001", "0110", "1101", "1100", "1100", "1101", "1110", "1101", "1010", "1110", "1100", "1001", "1011", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1111", "1110", "1110", "1111", "1111", "1111", "1111", "1111", "1111", "1111", "1110", "1110", "1110", "1110", "1110", "1111", "1010", "0100", "0101", "0011", "0010", "0010", "1001", "0110", "0001", "0001", "1001", "1101", "1011", "1001", "1100", "1001", "0110", "1011", "0111", "0100", "0111", "0110", "0101", "0111", "1000", "1001", "1001", "1000", "1100", "1011", "1010", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1110", "1110", "1110", "1111", "1111", "1111", "1110", "1011", "1011", "1100", "1111", "1111", "1110", "1111", "0111", "0011", "0101", "0100", "0011", "0010", "1010", "1110", "0110", "0001", "0101", "1101", "1100", "1100", "1011", "1001", "1010", "1001", "1001", "1001", "0110", "1000", "0111", "0101", "0011", "0011", "0011", "0010", "0101", "1011", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1110", "1110", "1110", "1110", "1111", "1111", "1110", "1110", "1101", "1111", "1111", "1111", "1111", "0101", "0100", "0011", "0100", "0011", "0010", "0011", "1000", "1100", "0111", "0100", "1001", "1101", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1010", "1001", "1000", "0110", "0101", "0101", "0011", "0011", "0100", "1100", "1101", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1111", "1110", "1111", "1111", "1111", "1111", "0101", "0010", "0010", "0010", "0011", "0011", "0100", "1001", "0110", "0101", "0001", "0010", "1010", "1101", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1010", "1001", "1000", "0110", "0100", "0100", "0001", "0101", "1100", "1101", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1111", "1111", "1111", "1111", "1111", "1111", "1000", "0000", "0000", "0001", "0001", "0010", "1001", "1001", "0011", "0101", "0010", "0110", "1010", "1010", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1011", "1010", "1010", "1001", "1000", "1000", "0111", "0110", "1101", "1110", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1100", "1000", "0010", "0001", "0001", "0001", "0110", "1100", "1010", "1000", "1010", "1101", "1101", "1100", "1011", "1010", "1011", "1100", "1100", "1011", "1011", "1011", "1011", "1010", "1010", "1001", "1001", "1000", "0111", "0111", "1010", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1011", "1010", "1100", "1010", "1011", "1110", "0110", "0000", "0001", "0011", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1011", "1010", "1001", "1100", "1100", "1011", "1011", "1011", "1011", "1010", "1001", "1001", "1000", "0111", "0111", "1100", "1100", "1100", "1100", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1011", "1011", "1101", "1011", "1011", "1011", "0000", "0001", "0001", "1000", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1011", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1010", "1010", "1100", "1100", "1100", "1100", "1101", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1100", "1100", "1101", "1001", "1001", "0010", "0000", "0000", "0001", "1011", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1100", "1101", "1101", "1100", "1100", "1011", "0100", "0000", "0001", "0010", "1000", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1100", "1110", "1110", "1100", "1100", "1000", "0010", "0011", "0011", "0011", "0111", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1101", "1110", "1110", "1101", "1100", "0111", "0011", "0001", "0101", "0010", "0111", "1101", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1110", "1101", "1101", "1110", "1101", "1101", "1110", "1110", "1110", "1101", "0110", "0010", "0100", "1000", "0100", "0100", "1001", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1011", "1100", "1101", "1101", "1101", "1110", "1110", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1110", "1110", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1110", "1101", "1110", "1010", "0110", "0001", "0100", "1000", "0111", "0010", "0100", "1010", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1110", "1110", "1110", "1110", "1101", "1101", "1101", "1101", "1110", "1100", "1101", "1110", "1101", "1101", "1001", "0110", "0010", "0010", "0110", "1001", "0101", "0001", "0110", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1101", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1101", "1110", "1110", "1110", "1101", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1110", "1100", "0111", "0110", "0011", "0001", "0101", "1011", "0111", "0010", "0110", "1011", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1110", "1101", "1110", "1110", "1101", "1101", "1101", "1110", "1110", "1110", "1110", "1110", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1101", "1101", "1101", "1001", "0111", "0111", "0100", "0000", "0011", "1001", "1001", "0110", "1011", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1110", "1101", "1101", "1101", "1110", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1000", "0111", "0111", "0100", "0100", "0100", "0111", "1011", "1011", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1011", "1101", "1101", "1101", "1100", "0111", "0111", "0111", "0110", "0100", "0100", "1011", "1011", "1011", "1100", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1110", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1101", "1101", "1101", "1010", "0111", "0111", "0111", "0101", "0100", "0110", "1000", "1011", "1100", "1100", "1101", "1101", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1011", "1101", "1101", "1101", "1101", "1001", "0111", "0111", "0111", "0111", "0111", "1001", "1000", "1011", "1101", "1100", "1100", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1011", "1100", "1100", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1011", "1101", "1101", "1101", "1100", "1000", "0111", "0111", "0111", "0111", "1000", "1010", "1000", "1011", "1101", "1100", "1100", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1101", "1101", "1101", "1011", "0111", "0111", "0111", "0111", "0111", "1000", "1001", "1000", "1011", "1101", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1100", "1101", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1011", "1100", "1101", "1101", "1101", "1001", "0111", "0111", "0111", "0111", "0111", "1000", "1010", "1010", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1011", "1101", "1101", "1101", "1100", "1000", "0111", "1000", "1000", "1000", "0111", "1000", "1010", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1011", "1011", "1011", "1011", "1011", "1011", "1011", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1101", "1101", "1100", "1100", "1100", "1100", "1100", "1101", "1100", "1100", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1101", "1100", "1100", "1101", "1101", "1101", "1011", "1000", "1000", "1000", "1000", "1000", "1000", "0111", "1001", "1100", "1100", "1100", "1100", "1100", "1100", "1100", "1100");
	

begin

	x <= conv_integer(x_control);
	y <= conv_integer(y_control);  


	process(clk,x,y)
	begin
		if clk'event and clk='1' then
			if (x < bredd + Xpos ) and (x > Xpos) and (y < hojd + Ypos) and (y > Ypos)  then
				counter <= (y-Ypos)*bredd + x - Xpos ; 
			end if;
			rgb_reg <= rgb_next;
		end if;
	end process;

	rgb_next <= ROM(counter) when (x < bredd + Xpos) and (x > Xpos )  and (y < hojd + Ypos) and (y > Ypos) else "1010";
	rgb<=rgb_reg;

	 
end Behavioral;
